library verilog;
use verilog.vl_types.all;
entity Block1_vlg_check_tst is
    port(
        y1              : in     vl_logic;
        y2              : in     vl_logic;
        y3              : in     vl_logic;
        y4              : in     vl_logic;
        y5              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Block1_vlg_check_tst;
