library verilog;
use verilog.vl_types.all;
entity Block1 is
    port(
        y1              : out    vl_logic;
        a               : in     vl_logic;
        b               : in     vl_logic;
        c               : in     vl_logic;
        y2              : out    vl_logic;
        d               : in     vl_logic;
        e               : in     vl_logic;
        y3              : out    vl_logic;
        f               : in     vl_logic;
        g               : in     vl_logic;
        y4              : out    vl_logic;
        h               : in     vl_logic;
        i               : in     vl_logic;
        y5              : out    vl_logic
    );
end Block1;
